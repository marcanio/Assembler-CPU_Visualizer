module ONES(ONE_OUTPUT);
output [15:0] ONE_OUTPUT;
assign ONE_OUTPUT[15:0]  = 16'b1111111111111111;

endmodule 