module BIOS_Hardcoded(b0,b1,b2,b3,b4,b5,b6,b7,b8,b9,b10,b11,b12,b13,b14,b15);

output [15:0] b0;
output [15:0] b1;
output [15:0] b2;
output [15:0] b3;
output [15:0] b4;
output [15:0] b5;
output [15:0] b6;
output [15:0] b7;
output [15:0] b8;
output [15:0] b9;
output [15:0] b10;
output [15:0] b11;
output [15:0] b12;
output [15:0] b13;
output [15:0] b14;
output [15:0] b15;

assign b0[15:0] = 16'b0000000000000000;
assign b1[15:0] = 16'b0000000000000000;
assign b2[15:0] = 16'b0000000000000000;
assign b3[15:0] = 16'b0000000000000000;
assign b4[15:0] = 16'b0000000000000000;
assign b5[15:0] = 16'b0000000000000000;
assign b6[15:0] = 16'b0000000000000000;
assign b7[15:0] = 16'b0000000000000000;
assign b8[15:0] = 16'b0000000000000000;
assign b9[15:0] = 16'b0000000000000000;
assign b10[15:0] = 16'b0000000000000000;
assign b11[15:0] = 16'b0000000000000000;
assign b12[15:0] = 16'b0000000000000000;
assign b13[15:0] = 16'b0000000000000000;
assign b14[15:0] = 16'b0000000000000000;
assign b15[15:0] = 16'b0000000000000000;

endmodule