module ZEROS(ZERO_OUTPUT);
output [7:0] ZERO_OUTPUT;
assign ZERO_OUTPUT[7:0]  = 8'b00000000;

endmodule 